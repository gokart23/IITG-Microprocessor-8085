----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    23:57:34 03/17/2015 
-- Design Name: 
-- Module Name:    ram - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.std_logic_arith.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity ram is
    Port ( cs : in  STD_LOGIC;
			  clk : in STD_LOGIC;
			  reset : in STD_LOGIC;
           en_read : in  STD_LOGIC;
           addr_bus : in  STD_LOGIC_VECTOR (15 downto 0);
           data_bus : inout  STD_LOGIC_VECTOR (7 downto 0));
end ram;

architecture ramArch of ram is
type ram_mem is array(0 to 127) of STD_LOGIC_VECTOR(7 downto 0);
signal ram : ram_mem;
begin
	process(reset, en_read, clk) begin
		if reset = '1' then
			-- load the ram with predef values
--			ram(256) <= "00000111";
--			ram(257) <= "00110001";
--			ram(258) <= "01000111";
--			ram(259) <= "00110010";
--			ram(260) <= "01001111";
--			ram(261) <= "00110011";
--			ram(262) <= "00100111";
--			ram(263) <= "00110100";
--			ram(264) <= "00001111";
--			ram(265) <= "11111111";
--			ram(512) <= x"02";
--			ram(513) <= x"02";
--			ram(514) <= x"03";
--			ram(515) <= x"04";
--			ram(516) <= x"05";
--ram(5) <= x"05";
--ram(10) <= "10000101";
--ram(11) <= "00000000";
--ram(12) <= "10000001";
--ram(13) <= "00000001";
--ram(14) <= "10000010";
--ram(15) <= "00000001";
--ram(16) <= "00000001";
--ram(17) <= "01010010";
--ram(18) <= "00001000";
--ram(19) <= "00000010";
--ram(20) <= "10100000";
--ram(21) <= "00000001";
--ram(22) <= "00010000";
--ram(23) <= "10000110";
--ram(24) <= "00000101";
--ram(25) <= "00011111";
--ram(26) <= "01001011";
--ram(27) <= "11011000";
--ram(28) <= "00000000";
--ram(29) <= "00010000";
--ram(30) <= "11001000";
--ram(31) <= "00000000";
--ram(32) <= "00010000";
--ram(33) <= "00000001";
--ram(34) <= "11111111";
--ram(10) <= "10000000";
--ram(11) <= "00000011";
--ram(12) <= "10000001";
--ram(13) <= "00001001";
--ram(14) <= "01000001";
--ram(15) <= "11111111";



--			ram(5) <= x"05";
--ram(10) <= "11000000";
--ram(11) <= "00000000";
--ram(12) <= "00110011";
--ram(13) <= "10000101";
--ram(14) <= "00000000";
--ram(15) <= "10000001";
--ram(16) <= "00000001";
--ram(17) <= "10000010";
--ram(18) <= "00000001";
--ram(19) <= "00000001";
--ram(20) <= "01010010";
--ram(21) <= "00001000";
--ram(22) <= "00000010";
--ram(23) <= "10100000";
--ram(24) <= "00000001";
--ram(25) <= "00010000";
--ram(26) <= "10000110";
--ram(27) <= "00000101";
--ram(28) <= "00011111";
--ram(29) <= "01001011";
--ram(30) <= "11011000";
--ram(31) <= "00000000";
--ram(32) <= "00010011";
--ram(33) <= "11001000";
--ram(34) <= "00000000";
--ram(35) <= "00010011";
--ram(36) <= "11101000";
--ram(37) <= "10000110";
--ram(38) <= "00110001";
--ram(39) <= "10000101";
--ram(40) <= "00000000";
--ram(41) <= "00111000";
--ram(42) <= "11101000";
--ram(43) <= "10000110";
--ram(44) <= "00110010";
--ram(45) <= "10000101";
--ram(46) <= "00000000";
--ram(47) <= "00111000";
--ram(48) <= "11000000";
--ram(49) <= "00000000";
--ram(50) <= "00000000";
--ram(51) <= "11100000";
--ram(52) <= "10000000";
--ram(53) <= "00111110";
--ram(54) <= "11100000";
--ram(55) <= "10000000";
--ram(56) <= "00000000";
--ram(57) <= "11100000";
--ram(58) <= "11000000";
--ram(59) <= "00000000";
--ram(60) <= "00001101";
--ram(61) <= "11101000";
--ram(62) <= "11111111";

--add em up
--ram(265) <= "00000101"; --earlier it was 508
--ram(261) <= "00000001";
--ram(260) <= "00000010";
--ram(259) <= "00000011";
--ram(258) <= "00000100";
--ram(257) <= "00000101";
--ram(256) <= "00000110";
--
--ram(8) <= "10000000";
--ram(9) <= "00000000";
--ram(10) <= "10000011";
--ram(11) <= "00000000";
--ram(12) <= "10000101";
--ram(13) <= "00000001";	
--ram(14) <= "10000110";
----ram(15) <= "11111100";
--ram(15) <= "00001001";
--ram(16) <= "00010111";
--ram(17) <= "00110010";
--ram(18) <= "00001111";
--ram(19) <= "00000011";
--ram(20) <= "01000001";
--ram(21) <= "00011000";
--ram(22) <= "00000010";
--ram(23) <= "10100100";
--ram(24) <= "00000001";
--ram(25) <= "00010000";
--ram(26) <= "11010000";
--ram(27) <= "00000000";
--ram(28) <= "00010001";
--ram(29) <= "00000011";
--ram(30) <= "11111111";

--alu test code
--ram(10) <= "10000001";
--ram(11) <= "00000101";
--ram(12) <= "10000000";
--ram(13) <= "00000011";
--ram(14) <= "01010001";
--ram(15) <= "01001001";
--ram(16) <= "11111111";

--fac with sub
ram(5) <= "00000101";
ram(10) <= "10000101";
ram(11) <= "00000000";
ram(12) <= "10000001";
ram(13) <= "00000001";
ram(14) <= "10000010";
ram(15) <= "00000001";
ram(16) <= "00000001";
ram(17) <= "01010010";
ram(18) <= "00001000";
ram(19) <= "00000010";
ram(20) <= "10100100";
ram(21) <= "11111111";
ram(22) <= "00010000";
ram(23) <= "10000110";
ram(24) <= "00000101";
ram(25) <= "00011111";
ram(26) <= "01001011";
ram(27) <= "11011000";
ram(28) <= "00000000";
ram(29) <= "00010000";
ram(30) <= "11001000";
ram(31) <= "00000000";
ram(32) <= "00010000";
ram(33) <= "00000001";
ram(34) <= "11111111";


----			ram(11) <= "10000000";
----			ram(12) <= "00000101";
----			ram(13) <= "10000001";
----			ram(14) <= "00000101";
----			ram(15) <= "01000001";
----			ram(16) <= "10100000";
----			ram(17) <= "00000101";
----			ram(18) <= "10000101";
----			ram(19) <= "00000000";
----			ram(20) <= "10000110";
----			ram(21) <= "00000101";
----			ram(22) <= "00111000";
--			ram(12) <= "00001111";
--			ram(13) <= "01000001";
--			ram(19) <= "11111111";
		elsif clk'event and clk = '1' and en_read = '1' and cs = '1' then 
			ram(conv_integer(unsigned(addr_bus))) <= data_bus;
		end if;
	end process;
	data_bus <= ram(conv_integer(unsigned(addr_bus))) when reset = '0' and en_read = '0' and cs = '1' else
					"ZZZZZZZZ";
end ramArch;

